// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Wed Jun 10 00:27:32 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [6:0] LEGUP_0 = 7'd0;
parameter [6:0] LEGUP_F_main_BB_entry_1 = 7'd1;
parameter [6:0] LEGUP_F_main_BB_while_body_i_2 = 7'd2;
parameter [6:0] LEGUP_F_main_BB_while_body_i_3 = 7'd3;
parameter [6:0] LEGUP_F_main_BB_while_body_i_4 = 7'd4;
parameter [6:0] LEGUP_F_main_BB_while_body_i16_preheader_5 = 7'd5;
parameter [6:0] LEGUP_F_main_BB_while_body_i16_6 = 7'd6;
parameter [6:0] LEGUP_F_main_BB_while_body_i16_7 = 7'd7;
parameter [6:0] LEGUP_F_main_BB_while_body_i16_8 = 7'd8;
parameter [6:0] LEGUP_F_main_BB_while_body_i10_preheader_9 = 7'd9;
parameter [6:0] LEGUP_F_main_BB_while_body_i10_10 = 7'd10;
parameter [6:0] LEGUP_F_main_BB_while_body_i10_11 = 7'd11;
parameter [6:0] LEGUP_F_main_BB_while_body_i4_preheader_12 = 7'd12;
parameter [6:0] LEGUP_F_main_BB_while_body_i4_13 = 7'd13;
parameter [6:0] LEGUP_F_main_BB_while_body_i4_14 = 7'd14;
parameter [6:0] LEGUP_F_main_BB_NodeBlock29_preheader_15 = 7'd15;
parameter [6:0] LEGUP_F_main_BB_NodeBlock29_16 = 7'd16;
parameter [6:0] LEGUP_F_main_BB_NodeBlock27_17 = 7'd17;
parameter [6:0] LEGUP_F_main_BB_NodeBlock25_18 = 7'd18;
parameter [6:0] LEGUP_F_main_BB_NodeBlock23_19 = 7'd19;
parameter [6:0] LEGUP_F_main_BB_LeafBlock21_20 = 7'd20;
parameter [6:0] LEGUP_F_main_BB_NodeBlock19_21 = 7'd21;
parameter [6:0] LEGUP_F_main_BB_NodeBlock17_22 = 7'd22;
parameter [6:0] LEGUP_F_main_BB_NodeBlock15_23 = 7'd23;
parameter [6:0] LEGUP_F_main_BB_NodeBlock13_24 = 7'd24;
parameter [6:0] LEGUP_F_main_BB_NodeBlock11_25 = 7'd25;
parameter [6:0] LEGUP_F_main_BB_NodeBlock9_26 = 7'd26;
parameter [6:0] LEGUP_F_main_BB_NodeBlock7_27 = 7'd27;
parameter [6:0] LEGUP_F_main_BB_NodeBlock5_28 = 7'd28;
parameter [6:0] LEGUP_F_main_BB_NodeBlock3_29 = 7'd29;
parameter [6:0] LEGUP_F_main_BB_NodeBlock1_30 = 7'd30;
parameter [6:0] LEGUP_F_main_BB_NodeBlock_31 = 7'd31;
parameter [6:0] LEGUP_F_main_BB_LeafBlock_32 = 7'd32;
parameter [6:0] LEGUP_F_main_BB_sw_bb1_33 = 7'd33;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_34 = 7'd34;
parameter [6:0] LEGUP_F_main_BB_if_else_35 = 7'd35;
parameter [6:0] LEGUP_F_main_BB_if_else_36 = 7'd36;
parameter [6:0] LEGUP_F_main_BB_sw_bb12_37 = 7'd37;
parameter [6:0] LEGUP_F_main_BB_if_else18_38 = 7'd38;
parameter [6:0] LEGUP_F_main_BB_if_else18_39 = 7'd39;
parameter [6:0] LEGUP_F_main_BB_sw_bb29_40 = 7'd40;
parameter [6:0] LEGUP_F_main_BB_sw_bb29_41 = 7'd41;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false_42 = 7'd42;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false_43 = 7'd43;
parameter [6:0] LEGUP_F_main_BB_sw_bb41_44 = 7'd44;
parameter [6:0] LEGUP_F_main_BB_sw_bb41_45 = 7'd45;
parameter [6:0] LEGUP_F_main_BB_if_then47_46 = 7'd46;
parameter [6:0] LEGUP_F_main_BB_if_then47_47 = 7'd47;
parameter [6:0] LEGUP_F_main_BB_if_then47_48 = 7'd48;
parameter [6:0] LEGUP_F_main_BB_if_end50_49 = 7'd49;
parameter [6:0] LEGUP_F_main_BB_if_end50_50 = 7'd50;
parameter [6:0] LEGUP_F_main_BB_sw_bb58_51 = 7'd51;
parameter [6:0] LEGUP_F_main_BB_sw_bb58_52 = 7'd52;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false64_53 = 7'd53;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false64_54 = 7'd54;
parameter [6:0] LEGUP_F_main_BB_sw_bb73_55 = 7'd55;
parameter [6:0] LEGUP_F_main_BB_sw_bb73_56 = 7'd56;
parameter [6:0] LEGUP_F_main_BB_if_then79_57 = 7'd57;
parameter [6:0] LEGUP_F_main_BB_if_then79_58 = 7'd58;
parameter [6:0] LEGUP_F_main_BB_if_then79_59 = 7'd59;
parameter [6:0] LEGUP_F_main_BB_if_end83_60 = 7'd60;
parameter [6:0] LEGUP_F_main_BB_if_end83_61 = 7'd61;
parameter [6:0] LEGUP_F_main_BB_sw_bb91_62 = 7'd62;
parameter [6:0] LEGUP_F_main_BB_if_else98_63 = 7'd63;
parameter [6:0] LEGUP_F_main_BB_if_else98_64 = 7'd64;
parameter [6:0] LEGUP_F_main_BB_sw_bb109_65 = 7'd65;
parameter [6:0] LEGUP_F_main_BB_sw_bb109_66 = 7'd66;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false115_67 = 7'd67;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false115_68 = 7'd68;
parameter [6:0] LEGUP_F_main_BB_sw_bb124_69 = 7'd69;
parameter [6:0] LEGUP_F_main_BB_sw_bb124_70 = 7'd70;
parameter [6:0] LEGUP_F_main_BB_if_then130_71 = 7'd71;
parameter [6:0] LEGUP_F_main_BB_if_then130_72 = 7'd72;
parameter [6:0] LEGUP_F_main_BB_if_then130_73 = 7'd73;
parameter [6:0] LEGUP_F_main_BB_if_end134_74 = 7'd74;
parameter [6:0] LEGUP_F_main_BB_if_end134_75 = 7'd75;
parameter [6:0] LEGUP_F_main_BB_sw_bb142_76 = 7'd76;
parameter [6:0] LEGUP_F_main_BB_sw_bb142_77 = 7'd77;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false148_78 = 7'd78;
parameter [6:0] LEGUP_F_main_BB_lor_lhs_false148_79 = 7'd79;
parameter [6:0] LEGUP_F_main_BB_sw_bb157_80 = 7'd80;
parameter [6:0] LEGUP_F_main_BB_sw_bb157_81 = 7'd81;
parameter [6:0] LEGUP_F_main_BB_if_then163_82 = 7'd82;
parameter [6:0] LEGUP_F_main_BB_if_then163_83 = 7'd83;
parameter [6:0] LEGUP_F_main_BB_if_then163_84 = 7'd84;
parameter [6:0] LEGUP_F_main_BB_if_end167_85 = 7'd85;
parameter [6:0] LEGUP_F_main_BB_if_end167_86 = 7'd86;
parameter [6:0] LEGUP_F_main_BB_sw_bb175_87 = 7'd87;
parameter [6:0] LEGUP_F_main_BB_sw_bb182_88 = 7'd88;
parameter [6:0] LEGUP_F_main_BB_sw_bb187_89 = 7'd89;
parameter [6:0] LEGUP_F_main_BB_sw_bb187_90 = 7'd90;
parameter [6:0] LEGUP_F_main_BB_sw_bb187_91 = 7'd91;
parameter [6:0] LEGUP_F_main_BB_sw_bb187_92 = 7'd92;
parameter [6:0] LEGUP_F_main_BB_if_else195_93 = 7'd93;
parameter [6:0] LEGUP_F_main_BB_if_else195_94 = 7'd94;
parameter [6:0] LEGUP_F_main_BB_if_else195_95 = 7'd95;
parameter [6:0] LEGUP_F_main_BB_sw_bb200_96 = 7'd96;
parameter [6:0] LEGUP_F_main_BB_NewDefault_97 = 7'd97;
parameter [6:0] LEGUP_F_main_BB_sw_epilog_98 = 7'd98;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [6:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [6:0] next_state;
wire  fsm_stall;
reg [6:0] main_while_body_i_indvar7;
reg [6:0] main_while_body_i_indvar7_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i_dt_04_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i_dt_04_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i_st_05_i;
reg [7:0] main_while_body_i_0;
reg [7:0] main_while_body_i_1;
reg [7:0] main_while_body_i_1_reg;
reg  main_while_body_i_exitcond;
reg  main_while_body_i_exitcond_reg;
reg [4:0] main_while_body_i16_indvar4;
reg [4:0] main_while_body_i16_indvar4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i16_dt_05_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i16_dt_05_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i16_st_06_i;
reg [31:0] main_while_body_i16_2;
reg [5:0] main_while_body_i16_3;
reg [5:0] main_while_body_i16_3_reg;
reg  main_while_body_i16_exitcond3;
reg  main_while_body_i16_exitcond3_reg;
reg [2:0] main_while_body_i10_indvar1;
reg [2:0] main_while_body_i10_indvar1_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i10_s_010_i5;
reg [3:0] main_while_body_i10_4;
reg [3:0] main_while_body_i10_4_reg;
reg  main_while_body_i10_exitcond2;
reg  main_while_body_i10_exitcond2_reg;
reg [2:0] main_while_body_i4_indvar;
reg [2:0] main_while_body_i4_indvar_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_while_body_i4_s_010_i;
reg [3:0] main_while_body_i4_5;
reg [3:0] main_while_body_i4_5_reg;
reg  main_while_body_i4_exitcond1;
reg  main_while_body_i4_exitcond1_reg;
reg [31:0] main_NodeBlock29_state_0;
reg [31:0] main_NodeBlock29_state_0_reg;
reg [31:0] main_NodeBlock29_current_sroa_30_0;
reg [31:0] main_NodeBlock29_current_sroa_30_0_reg;
reg [31:0] main_NodeBlock29_current_sroa_0_0;
reg [31:0] main_NodeBlock29_current_sroa_0_0_reg;
reg [31:0] main_NodeBlock29_inputIndex_0;
reg [31:0] main_NodeBlock29_inputIndex_0_reg;
reg [31:0] main_NodeBlock29_stackIndex_0;
reg [31:0] main_NodeBlock29_stackIndex_0_reg;
reg  main_NodeBlock29_modified_0;
reg  main_NodeBlock29_modified_0_reg;
reg  main_NodeBlock29_firstEdge_0;
reg  main_NodeBlock29_firstEdge_0_reg;
reg [31:0] main_NodeBlock29_next_state_0;
reg [31:0] main_NodeBlock29_next_state_0_reg;
reg [7:0] main_NodeBlock29_next_modified_0;
reg [7:0] main_NodeBlock29_next_modified_0_reg;
reg [7:0] main_NodeBlock29_next_firstEdge_0;
reg [7:0] main_NodeBlock29_next_firstEdge_0_reg;
reg [1:0] main_NodeBlock29_bit_select15;
reg [1:0] main_NodeBlock29_bit_select15_reg;
reg [1:0] main_NodeBlock29_bit_select13;
reg [1:0] main_NodeBlock29_bit_select13_reg;
reg [29:0] main_NodeBlock29_bit_select11;
reg [29:0] main_NodeBlock29_bit_select11_reg;
reg [29:0] main_NodeBlock29_bit_select9;
reg [29:0] main_NodeBlock29_bit_select9_reg;
reg [29:0] main_NodeBlock29_bit_select5;
reg [29:0] main_NodeBlock29_bit_select5_reg;
reg  main_NodeBlock29_Pivot30;
reg  main_NodeBlock27_Pivot28;
reg  main_NodeBlock25_Pivot26;
reg  main_NodeBlock23_Pivot24;
reg  main_LeafBlock21_SwitchLeaf22;
reg  main_NodeBlock19_Pivot20;
reg  main_NodeBlock17_Pivot18;
reg  main_NodeBlock15_Pivot16;
reg [31:0] main_NodeBlock15_bit_concat23;
reg [31:0] main_NodeBlock15_bit_concat23_reg;
reg  main_NodeBlock13_Pivot14;
reg  main_NodeBlock11_Pivot12;
reg  main_NodeBlock9_Pivot10;
reg  main_NodeBlock7_Pivot8;
reg [31:0] main_NodeBlock7_bit_concat22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_NodeBlock7_arrayidx32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_NodeBlock7_arrayidx32_reg;
reg  main_NodeBlock5_Pivot6;
reg [31:0] main_NodeBlock5_bit_concat21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_NodeBlock5_arrayidx62;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_NodeBlock5_arrayidx62_reg;
reg  main_NodeBlock3_Pivot4;
reg  main_NodeBlock1_Pivot2;
reg  main_NodeBlock_Pivot;
reg  main_LeafBlock_SwitchLeaf;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb1_arrayidx;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb1_arrayidx_reg;
reg [15:0] main_sw_bb1_6;
reg  main_sw_bb1_bit_select19;
reg [31:0] main_sw_bb1_bit_concat20;
reg  main_sw_bb1_cmp;
reg [31:0] main_sw_bb1_add8_pre;
reg [31:0] main_sw_bb1_add8_pre_reg;
reg [15:0] main_land_lhs_true_7;
reg  main_land_lhs_true_bit_select17;
reg [31:0] main_land_lhs_true_bit_concat18;
reg  main_land_lhs_true_cmp4;
reg [31:0] main_if_else_8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_else_arrayidx9;
reg [31:0] main_if_else_9;
reg [31:0] main_if_else_add11;
reg [31:0] main_if_else_add11_reg;
reg [31:0] main_sw_bb12_bit_concat16;
reg [31:0] main_sw_bb12_bit_concat16_reg;
reg [31:0] main_sw_bb12_bit_concat14;
reg [31:0] main_sw_bb12_bit_concat14_reg;
reg  main_sw_bb12_cmp16;
reg [31:0] main_if_else18_sub;
reg  main_if_else18_cmp24;
reg  main_if_else18_cmp24_reg;
reg [2:0] main_if_else18_1;
reg [7:0] main_sw_bb29_10;
reg  main_sw_bb29_tobool;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_lor_lhs_false_arrayidx34;
reg [31:0] main_lor_lhs_false_11;
reg  main_lor_lhs_false_cmp35_not;
reg  main_lor_lhs_false_brmerge;
reg [3:0] main_lor_lhs_false_292;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then47_arrayidx49;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then47_arrayidx49_reg;
reg [31:0] main_if_then47_12;
reg [31:0] main_if_then47_inc;
reg [31:0] main_if_end50_add52;
reg [31:0] main_if_end50_add52_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end50_arrayidx55;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end50_arrayidx56;
reg [31:0] main_if_end50_add57;
reg [31:0] main_if_end50_add57_reg;
reg [7:0] main_sw_bb58_13;
reg  main_sw_bb58_tobool63;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_lor_lhs_false64_arrayidx66;
reg [31:0] main_lor_lhs_false64_14;
reg  main_lor_lhs_false64_cmp67_not;
reg  main_lor_lhs_false64_brmerge286;
reg [3:0] main_lor_lhs_false64_293;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then79_arrayidx81;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then79_arrayidx81_reg;
reg [31:0] main_if_then79_15;
reg [31:0] main_if_then79_inc82;
reg [31:0] main_if_end83_sub85;
reg [31:0] main_if_end83_sub85_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end83_arrayidx88;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end83_arrayidx89;
reg [31:0] main_if_end83_add90;
reg [31:0] main_if_end83_add90_reg;
reg [31:0] main_sw_bb91_bit_concat12;
reg [31:0] main_sw_bb91_bit_concat12_reg;
reg [31:0] main_sw_bb91_bit_concat10;
reg [31:0] main_sw_bb91_bit_concat10_reg;
reg  main_sw_bb91_cmp96;
reg [31:0] main_if_else98_sub95;
reg  main_if_else98_cmp104;
reg  main_if_else98_cmp104_reg;
reg [3:0] main_if_else98_287;
reg [31:0] main_sw_bb109_bit_concat8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb109_arrayidx113;
reg [7:0] main_sw_bb109_16;
reg  main_sw_bb109_tobool114;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_lor_lhs_false115_arrayidx117;
reg [31:0] main_lor_lhs_false115_17;
reg  main_lor_lhs_false115_cmp118_not;
reg  main_lor_lhs_false115_brmerge288;
reg [3:0] main_lor_lhs_false115_294;
reg [31:0] main_sw_bb124_bit_concat7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb124_arrayidx128;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then130_arrayidx132;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then130_arrayidx132_reg;
reg [31:0] main_if_then130_18;
reg [31:0] main_if_then130_inc133;
reg [31:0] main_if_end134_add136;
reg [31:0] main_if_end134_add136_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end134_arrayidx139;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end134_arrayidx140;
reg [31:0] main_if_end134_add141;
reg [31:0] main_if_end134_add141_reg;
reg [31:0] main_sw_bb142_bit_concat6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb142_arrayidx146;
reg [7:0] main_sw_bb142_19;
reg  main_sw_bb142_tobool147;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_lor_lhs_false148_arrayidx150;
reg [31:0] main_lor_lhs_false148_20;
reg  main_lor_lhs_false148_cmp151_not;
reg  main_lor_lhs_false148_brmerge289;
reg [3:0] main_lor_lhs_false148_295;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb157_arrayidx161;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then163_arrayidx165;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then163_arrayidx165_reg;
reg [31:0] main_if_then163_21;
reg [31:0] main_if_then163_inc166;
reg [31:0] main_if_end167_sub169;
reg [31:0] main_if_end167_sub169_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end167_arrayidx172;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end167_arrayidx173;
reg [31:0] main_if_end167_add174;
reg [31:0] main_if_end167_add174_reg;
reg  main_sw_bb175_cmp178;
reg [3:0] main_sw_bb175_290;
reg [3:0] main_sw_bb182_291;
reg [7:0] main_sw_bb182_next_modified_0;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb187_arrayidx188;
reg [31:0] main_sw_bb187_22;
reg [31:0] main_sw_bb187_22_reg;
reg [29:0] main_sw_bb187_bit_select3;
reg [31:0] main_sw_bb187_bit_concat4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb187_arrayidx190;
reg [31:0] main_sw_bb187_23;
reg [31:0] main_sw_bb187_add191;
reg [31:0] main_sw_bb187_add191_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_sw_bb187_arrayidx192;
reg  main_sw_bb187_cmp193;
reg  main_sw_bb187_cmp193_reg;
reg [31:0] main_if_else195_sub196;
reg [31:0] main_if_else195_sub196_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_else195_arrayidx198;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_else195_arrayidx198_reg;
reg [31:0] main_if_else195_24;
reg [31:0] main_if_else195_dec;
reg [31:0] main_sw_epilog_next_state_1;
reg [31:0] main_sw_epilog_next_state_1_reg;
reg [31:0] main_sw_epilog_next_current_sroa_6_1;
reg [31:0] main_sw_epilog_next_current_sroa_6_1_reg;
reg [31:0] main_sw_epilog_next_current_sroa_0_1;
reg [31:0] main_sw_epilog_next_current_sroa_0_1_reg;
reg [31:0] main_sw_epilog_next_inputIndex_1;
reg [31:0] main_sw_epilog_next_inputIndex_1_reg;
reg [31:0] main_sw_epilog_next_stackIndex_1;
reg [31:0] main_sw_epilog_next_stackIndex_1_reg;
reg [7:0] main_sw_epilog_next_modified_1;
reg [7:0] main_sw_epilog_next_modified_1_reg;
reg [7:0] main_sw_epilog_next_firstEdge_1;
reg [7:0] main_sw_epilog_next_firstEdge_1_reg;
reg  main_sw_epilog_bit_select1;
reg  main_sw_epilog_bit_select;
reg [7:0] main_sw_epilog_bit_concat2;
reg  main_sw_epilog_phitmp;
reg [7:0] main_sw_epilog_bit_concat;
reg  main_sw_epilog_phitmp279;
reg [3:0] main_input_address_a;
wire [31:0] main_input_out_a;
reg [3:0] main_input_address_b;
wire [31:0] main_input_out_b;
reg [5:0] main_grid_address_a;
wire [7:0] main_grid_out_a;
wire [5:0] main_grid_address_b;
wire [7:0] main_grid_out_b;
reg [3:0] main_bypass_address_a;
wire [31:0] main_bypass_out_a;
wire [3:0] main_bypass_address_b;
wire [31:0] main_bypass_out_b;
reg [5:0] main_entry_grid_address_a;
reg  main_entry_grid_write_enable_a;
reg [7:0] main_entry_grid_in_a;
wire [7:0] main_entry_grid_out_a;
reg [3:0] main_entry_bypass_address_a;
reg  main_entry_bypass_write_enable_a;
reg [31:0] main_entry_bypass_in_a;
wire [31:0] main_entry_bypass_out_a;
reg [2:0] main_entry_stackNode_address_a;
reg  main_entry_stackNode_write_enable_a;
reg [31:0] main_entry_stackNode_in_a;
wire [31:0] main_entry_stackNode_out_a;
reg [2:0] main_entry_stackOutput_address_a;
reg  main_entry_stackOutput_write_enable_a;
reg [31:0] main_entry_stackOutput_in_a;
wire [31:0] main_entry_stackOutput_out_a;
wire [5:0] main_NodeBlock29_Pivot30_op1_temp;
wire [5:0] main_NodeBlock27_Pivot28_op1_temp;
wire [5:0] main_NodeBlock25_Pivot26_op1_temp;
wire [5:0] main_NodeBlock23_Pivot24_op1_temp;
wire [5:0] main_NodeBlock19_Pivot20_op1_temp;
wire [5:0] main_NodeBlock17_Pivot18_op1_temp;
wire [5:0] main_NodeBlock15_Pivot16_op1_temp;
wire [1:0] main_NodeBlock15_bit_concat23_bit_select_operand_2;
wire [5:0] main_NodeBlock13_Pivot14_op1_temp;
wire [4:0] main_NodeBlock11_Pivot12_op1_temp;
wire [4:0] main_NodeBlock9_Pivot10_op1_temp;
wire [4:0] main_NodeBlock7_Pivot8_op1_temp;
wire [1:0] main_NodeBlock7_bit_concat22_bit_select_operand_2;
wire [4:0] main_NodeBlock5_Pivot6_op1_temp;
wire [1:0] main_NodeBlock5_bit_concat21_bit_select_operand_2;
wire [3:0] main_NodeBlock3_Pivot4_op1_temp;
wire [3:0] main_NodeBlock1_Pivot2_op1_temp;
wire [2:0] main_NodeBlock_Pivot_op1_temp;
wire [30:0] main_sw_bb1_bit_concat20_bit_select_operand_0;
wire [30:0] main_land_lhs_true_bit_concat18_bit_select_operand_0;
wire [29:0] main_sw_bb12_bit_concat16_bit_select_operand_0;
wire [29:0] main_sw_bb12_bit_concat14_bit_select_operand_0;
wire [1:0] main_if_else18_cmp24_op1_temp;
wire [1:0] main_sw_bb91_bit_concat12_bit_select_operand_0;
wire [1:0] main_sw_bb91_bit_concat10_bit_select_operand_0;
wire [1:0] main_if_else98_cmp104_op1_temp;
wire [1:0] main_sw_bb109_bit_concat8_bit_select_operand_2;
wire [1:0] main_sw_bb124_bit_concat7_bit_select_operand_2;
wire [1:0] main_sw_bb142_bit_concat6_bit_select_operand_2;
wire [1:0] main_sw_bb187_bit_concat4_bit_select_operand_2;
wire [6:0] main_sw_epilog_bit_concat2_bit_select_operand_0;
wire [6:0] main_sw_epilog_bit_concat_bit_select_operand_0;



// @main.input = private unnamed_addr constant [16 x i32] [i32 0, i32 2, i32 0, i32 8, i32 2, i32 2, i32 1, i32 9, i32 9, i32 2, i32 6, i32 11, i32 11, i32 2, i32 0, i32 0], align 4
rom_dual_port main_input (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_input_address_a ),
	.q_a( main_input_out_a ),
	.address_b( main_input_address_b ),
	.q_b( main_input_out_b )
);
defparam main_input.width_a = 32;
defparam main_input.widthad_a = 4;
defparam main_input.numwords_a = 16;
defparam main_input.width_b = 32;
defparam main_input.widthad_b = 4;
defparam main_input.numwords_b = 16;
defparam main_input.latency = 1;
defparam main_input.init_file = {`MEM_INIT_DIR, "main_input.mif"};


// @main.grid = private unnamed_addr constant [64 x i8] c"\00\00\00\00\00\00\00\00\00\00\00\01\00\00\00\00\01\00\00\01\01\00\00\01\00\00\00\00\00\00\00\00\00\00\00\00\00\00\00\01\00\00\00\00\00\01\00\00\...
rom_dual_port main_grid (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_grid_address_a ),
	.q_a( main_grid_out_a ),
	.address_b( main_grid_address_b ),
	.q_b( main_grid_out_b )
);
defparam main_grid.width_a = 8;
defparam main_grid.widthad_a = 6;
defparam main_grid.numwords_a = 64;
defparam main_grid.width_b = 8;
defparam main_grid.widthad_b = 6;
defparam main_grid.numwords_b = 64;
defparam main_grid.latency = 1;
defparam main_grid.init_file = {`MEM_INIT_DIR, "main_grid.mif"};


// @main.bypass = private unnamed_addr constant [16 x i32] [i32 1, i32 1, i32 1, i32 1, i32 1, i32 1, i32 1, i32 0, i32 1, i32 1, i32 1, i32 1, i32 0, i32 1, i32 0, i32 1], align 4
rom_dual_port main_bypass (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_bypass_address_a ),
	.q_a( main_bypass_out_a ),
	.address_b( main_bypass_address_b ),
	.q_b( main_bypass_out_b )
);
defparam main_bypass.width_a = 32;
defparam main_bypass.widthad_a = 4;
defparam main_bypass.numwords_a = 16;
defparam main_bypass.width_b = 32;
defparam main_bypass.widthad_b = 4;
defparam main_bypass.numwords_b = 16;
defparam main_bypass.latency = 1;
defparam main_bypass.init_file = {`MEM_INIT_DIR, "main_bypass.mif"};


//   %grid = alloca [64 x i8], align 1, !MSB !46, !LSB !47, !extendFrom !46
ram_single_port_intel main_entry_grid (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_grid_address_a ),
	.wren_a( main_entry_grid_write_enable_a ),
	.data_a( main_entry_grid_in_a ),
	.byteena_a( {1{1'b1}} ),
	.q_a( main_entry_grid_out_a )
);
defparam main_entry_grid.width_a = 8;
defparam main_entry_grid.widthad_a = 6;
defparam main_entry_grid.width_be_a = 1;
defparam main_entry_grid.numwords_a = 64;
defparam main_entry_grid.latency = 1;


//   %bypass = alloca [16 x i32], align 4, !MSB !46, !LSB !47, !extendFrom !46
ram_single_port_intel main_entry_bypass (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_bypass_address_a ),
	.wren_a( main_entry_bypass_write_enable_a ),
	.data_a( main_entry_bypass_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_bypass_out_a )
);
defparam main_entry_bypass.width_a = 32;
defparam main_entry_bypass.widthad_a = 4;
defparam main_entry_bypass.width_be_a = 4;
defparam main_entry_bypass.numwords_a = 16;
defparam main_entry_bypass.latency = 1;


//   %stackNode = alloca [6 x i32], align 4, !MSB !46, !LSB !47, !extendFrom !46
ram_single_port_intel main_entry_stackNode (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_stackNode_address_a ),
	.wren_a( main_entry_stackNode_write_enable_a ),
	.data_a( main_entry_stackNode_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_stackNode_out_a )
);
defparam main_entry_stackNode.width_a = 32;
defparam main_entry_stackNode.widthad_a = 3;
defparam main_entry_stackNode.width_be_a = 4;
defparam main_entry_stackNode.numwords_a = 6;
defparam main_entry_stackNode.latency = 1;


//   %stackOutput = alloca [6 x i32], align 4, !MSB !46, !LSB !47, !extendFrom !46
ram_single_port_intel main_entry_stackOutput (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_stackOutput_address_a ),
	.wren_a( main_entry_stackOutput_write_enable_a ),
	.data_a( main_entry_stackOutput_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_stackOutput_out_a )
);
defparam main_entry_stackOutput.width_a = 32;
defparam main_entry_stackOutput.widthad_a = 3;
defparam main_entry_stackOutput.width_be_a = 4;
defparam main_entry_stackOutput.numwords_a = 6;
defparam main_entry_stackOutput.latency = 1;

always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_LeafBlock21_20:
	if ((fsm_stall == 1'd0) && (main_LeafBlock21_SwitchLeaf22 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb187_89;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock21_SwitchLeaf22 == 1'd0))
		next_state = LEGUP_F_main_BB_NewDefault_97;
LEGUP_F_main_BB_LeafBlock_32:
	if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd1))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd0))
		next_state = LEGUP_F_main_BB_NewDefault_97;
LEGUP_F_main_BB_NewDefault_97:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_NodeBlock11_25:
	if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock3_29;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock9_26;
LEGUP_F_main_BB_NodeBlock13_24:
	if ((fsm_stall == 1'd0) && (main_NodeBlock13_Pivot14 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb91_62;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock13_Pivot14 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb142_76;
LEGUP_F_main_BB_NodeBlock15_23:
	if ((fsm_stall == 1'd0) && (main_NodeBlock15_Pivot16 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb157_80;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock15_Pivot16 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb109_65;
LEGUP_F_main_BB_NodeBlock17_22:
	if ((fsm_stall == 1'd0) && (main_NodeBlock17_Pivot18 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock13_24;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock17_Pivot18 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock15_23;
LEGUP_F_main_BB_NodeBlock19_21:
	if ((fsm_stall == 1'd0) && (main_NodeBlock19_Pivot20 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb124_69;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock19_Pivot20 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb175_87;
LEGUP_F_main_BB_NodeBlock1_30:
	if ((fsm_stall == 1'd0) && (main_NodeBlock1_Pivot2 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb200_96;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock1_Pivot2 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb12_37;
LEGUP_F_main_BB_NodeBlock23_19:
	if ((fsm_stall == 1'd0) && (main_NodeBlock23_Pivot24 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb182_88;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock23_Pivot24 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock21_20;
LEGUP_F_main_BB_NodeBlock25_18:
	if ((fsm_stall == 1'd0) && (main_NodeBlock25_Pivot26 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock19_21;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock25_Pivot26 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock23_19;
LEGUP_F_main_BB_NodeBlock27_17:
	if ((fsm_stall == 1'd0) && (main_NodeBlock27_Pivot28 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock17_22;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock27_Pivot28 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock25_18;
LEGUP_F_main_BB_NodeBlock29_16:
	if ((fsm_stall == 1'd0) && (main_NodeBlock29_Pivot30 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock11_25;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock29_Pivot30 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock27_17;
LEGUP_F_main_BB_NodeBlock29_preheader_15:
		next_state = LEGUP_F_main_BB_NodeBlock29_16;
LEGUP_F_main_BB_NodeBlock3_29:
	if ((fsm_stall == 1'd0) && (main_NodeBlock3_Pivot4 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock_31;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock3_Pivot4 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock1_30;
LEGUP_F_main_BB_NodeBlock5_28:
	if ((fsm_stall == 1'd0) && (main_NodeBlock5_Pivot6 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb58_51;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock5_Pivot6 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb73_55;
LEGUP_F_main_BB_NodeBlock7_27:
	if ((fsm_stall == 1'd0) && (main_NodeBlock7_Pivot8 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_bb29_40;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock7_Pivot8 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb41_44;
LEGUP_F_main_BB_NodeBlock9_26:
	if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock5_28;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock7_27;
LEGUP_F_main_BB_NodeBlock_31:
	if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock_32;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd0))
		next_state = LEGUP_F_main_BB_sw_bb1_33;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_while_body_i_2;
LEGUP_F_main_BB_if_else18_38:
		next_state = LEGUP_F_main_BB_if_else18_39;
LEGUP_F_main_BB_if_else18_39:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_else195_93:
		next_state = LEGUP_F_main_BB_if_else195_94;
LEGUP_F_main_BB_if_else195_94:
		next_state = LEGUP_F_main_BB_if_else195_95;
LEGUP_F_main_BB_if_else195_95:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_else98_63:
		next_state = LEGUP_F_main_BB_if_else98_64;
LEGUP_F_main_BB_if_else98_64:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_else_35:
		next_state = LEGUP_F_main_BB_if_else_36;
LEGUP_F_main_BB_if_else_36:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_end134_74:
		next_state = LEGUP_F_main_BB_if_end134_75;
LEGUP_F_main_BB_if_end134_75:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_end167_85:
		next_state = LEGUP_F_main_BB_if_end167_86;
LEGUP_F_main_BB_if_end167_86:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_end50_49:
		next_state = LEGUP_F_main_BB_if_end50_50;
LEGUP_F_main_BB_if_end50_50:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_end83_60:
		next_state = LEGUP_F_main_BB_if_end83_61;
LEGUP_F_main_BB_if_end83_61:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_if_then130_71:
		next_state = LEGUP_F_main_BB_if_then130_72;
LEGUP_F_main_BB_if_then130_72:
		next_state = LEGUP_F_main_BB_if_then130_73;
LEGUP_F_main_BB_if_then130_73:
		next_state = LEGUP_F_main_BB_if_end134_74;
LEGUP_F_main_BB_if_then163_82:
		next_state = LEGUP_F_main_BB_if_then163_83;
LEGUP_F_main_BB_if_then163_83:
		next_state = LEGUP_F_main_BB_if_then163_84;
LEGUP_F_main_BB_if_then163_84:
		next_state = LEGUP_F_main_BB_if_end167_85;
LEGUP_F_main_BB_if_then47_46:
		next_state = LEGUP_F_main_BB_if_then47_47;
LEGUP_F_main_BB_if_then47_47:
		next_state = LEGUP_F_main_BB_if_then47_48;
LEGUP_F_main_BB_if_then47_48:
		next_state = LEGUP_F_main_BB_if_end50_49;
LEGUP_F_main_BB_if_then79_57:
		next_state = LEGUP_F_main_BB_if_then79_58;
LEGUP_F_main_BB_if_then79_58:
		next_state = LEGUP_F_main_BB_if_then79_59;
LEGUP_F_main_BB_if_then79_59:
		next_state = LEGUP_F_main_BB_if_end83_60;
LEGUP_F_main_BB_land_lhs_true_34:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true_cmp4 == 1'd1))
		next_state = LEGUP_F_main_BB_if_else_35;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true_cmp4 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_lor_lhs_false115_67:
		next_state = LEGUP_F_main_BB_lor_lhs_false115_68;
LEGUP_F_main_BB_lor_lhs_false115_68:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_lor_lhs_false148_78:
		next_state = LEGUP_F_main_BB_lor_lhs_false148_79;
LEGUP_F_main_BB_lor_lhs_false148_79:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_lor_lhs_false64_53:
		next_state = LEGUP_F_main_BB_lor_lhs_false64_54;
LEGUP_F_main_BB_lor_lhs_false64_54:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_lor_lhs_false_42:
		next_state = LEGUP_F_main_BB_lor_lhs_false_43;
LEGUP_F_main_BB_lor_lhs_false_43:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb109_65:
		next_state = LEGUP_F_main_BB_sw_bb109_66;
LEGUP_F_main_BB_sw_bb109_66:
	if ((fsm_stall == 1'd0) && (main_sw_bb109_tobool114 == 1'd1))
		next_state = LEGUP_F_main_BB_lor_lhs_false115_67;
	else if ((fsm_stall == 1'd0) && (main_sw_bb109_tobool114 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb124_69:
		next_state = LEGUP_F_main_BB_sw_bb124_70;
LEGUP_F_main_BB_sw_bb124_70:
	if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_end134_74;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_then130_71;
LEGUP_F_main_BB_sw_bb12_37:
	if ((fsm_stall == 1'd0) && (main_sw_bb12_cmp16 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
	else if ((fsm_stall == 1'd0) && (main_sw_bb12_cmp16 == 1'd0))
		next_state = LEGUP_F_main_BB_if_else18_38;
LEGUP_F_main_BB_sw_bb142_76:
		next_state = LEGUP_F_main_BB_sw_bb142_77;
LEGUP_F_main_BB_sw_bb142_77:
	if ((fsm_stall == 1'd0) && (main_sw_bb142_tobool147 == 1'd1))
		next_state = LEGUP_F_main_BB_lor_lhs_false148_78;
	else if ((fsm_stall == 1'd0) && (main_sw_bb142_tobool147 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb157_80:
		next_state = LEGUP_F_main_BB_sw_bb157_81;
LEGUP_F_main_BB_sw_bb157_81:
	if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_end167_85;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_then163_82;
LEGUP_F_main_BB_sw_bb175_87:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb182_88:
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb187_89:
		next_state = LEGUP_F_main_BB_sw_bb187_90;
LEGUP_F_main_BB_sw_bb187_90:
		next_state = LEGUP_F_main_BB_sw_bb187_91;
LEGUP_F_main_BB_sw_bb187_91:
		next_state = LEGUP_F_main_BB_sw_bb187_92;
LEGUP_F_main_BB_sw_bb187_92:
	if ((fsm_stall == 1'd0) && (main_sw_bb187_cmp193_reg == 1'd1))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
	else if ((fsm_stall == 1'd0) && (main_sw_bb187_cmp193_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_else195_93;
LEGUP_F_main_BB_sw_bb1_33:
	if ((fsm_stall == 1'd0) && (main_sw_bb1_cmp == 1'd1))
		next_state = LEGUP_F_main_BB_if_else_35;
	else if ((fsm_stall == 1'd0) && (main_sw_bb1_cmp == 1'd0))
		next_state = LEGUP_F_main_BB_land_lhs_true_34;
LEGUP_F_main_BB_sw_bb200_96:
		next_state = LEGUP_0;
LEGUP_F_main_BB_sw_bb29_40:
		next_state = LEGUP_F_main_BB_sw_bb29_41;
LEGUP_F_main_BB_sw_bb29_41:
	if ((fsm_stall == 1'd0) && (main_sw_bb29_tobool == 1'd1))
		next_state = LEGUP_F_main_BB_lor_lhs_false_42;
	else if ((fsm_stall == 1'd0) && (main_sw_bb29_tobool == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb41_44:
		next_state = LEGUP_F_main_BB_sw_bb41_45;
LEGUP_F_main_BB_sw_bb41_45:
	if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_end50_49;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_then47_46;
LEGUP_F_main_BB_sw_bb58_51:
		next_state = LEGUP_F_main_BB_sw_bb58_52;
LEGUP_F_main_BB_sw_bb58_52:
	if ((fsm_stall == 1'd0) && (main_sw_bb58_tobool63 == 1'd1))
		next_state = LEGUP_F_main_BB_lor_lhs_false64_53;
	else if ((fsm_stall == 1'd0) && (main_sw_bb58_tobool63 == 1'd0))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
LEGUP_F_main_BB_sw_bb73_55:
		next_state = LEGUP_F_main_BB_sw_bb73_56;
LEGUP_F_main_BB_sw_bb73_56:
	if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_end83_60;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock29_firstEdge_0_reg == 1'd0))
		next_state = LEGUP_F_main_BB_if_then79_57;
LEGUP_F_main_BB_sw_bb91_62:
	if ((fsm_stall == 1'd0) && (main_sw_bb91_cmp96 == 1'd1))
		next_state = LEGUP_F_main_BB_sw_epilog_98;
	else if ((fsm_stall == 1'd0) && (main_sw_bb91_cmp96 == 1'd0))
		next_state = LEGUP_F_main_BB_if_else98_63;
LEGUP_F_main_BB_sw_epilog_98:
		next_state = LEGUP_F_main_BB_NodeBlock29_16;
LEGUP_F_main_BB_while_body_i10_10:
		next_state = LEGUP_F_main_BB_while_body_i10_11;
LEGUP_F_main_BB_while_body_i10_11:
	if ((fsm_stall == 1'd0) && (main_while_body_i10_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_while_body_i4_preheader_12;
	else if ((fsm_stall == 1'd0) && (main_while_body_i10_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i10_10;
LEGUP_F_main_BB_while_body_i10_preheader_9:
		next_state = LEGUP_F_main_BB_while_body_i10_10;
LEGUP_F_main_BB_while_body_i16_6:
		next_state = LEGUP_F_main_BB_while_body_i16_7;
LEGUP_F_main_BB_while_body_i16_7:
		next_state = LEGUP_F_main_BB_while_body_i16_8;
LEGUP_F_main_BB_while_body_i16_8:
	if ((fsm_stall == 1'd0) && (main_while_body_i16_exitcond3_reg == 1'd1))
		next_state = LEGUP_F_main_BB_while_body_i10_preheader_9;
	else if ((fsm_stall == 1'd0) && (main_while_body_i16_exitcond3_reg == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i16_6;
LEGUP_F_main_BB_while_body_i16_preheader_5:
		next_state = LEGUP_F_main_BB_while_body_i16_6;
LEGUP_F_main_BB_while_body_i4_13:
		next_state = LEGUP_F_main_BB_while_body_i4_14;
LEGUP_F_main_BB_while_body_i4_14:
	if ((fsm_stall == 1'd0) && (main_while_body_i4_exitcond1_reg == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock29_preheader_15;
	else if ((fsm_stall == 1'd0) && (main_while_body_i4_exitcond1_reg == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i4_13;
LEGUP_F_main_BB_while_body_i4_preheader_12:
		next_state = LEGUP_F_main_BB_while_body_i4_13;
LEGUP_F_main_BB_while_body_i_2:
		next_state = LEGUP_F_main_BB_while_body_i_3;
LEGUP_F_main_BB_while_body_i_3:
		next_state = LEGUP_F_main_BB_while_body_i_4;
LEGUP_F_main_BB_while_body_i_4:
	if ((fsm_stall == 1'd0) && (main_while_body_i_exitcond_reg == 1'd1))
		next_state = LEGUP_F_main_BB_while_body_i16_preheader_5;
	else if ((fsm_stall == 1'd0) && (main_while_body_i_exitcond_reg == 1'd0))
		next_state = LEGUP_F_main_BB_while_body_i_2;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar7 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_body_i_4) & (fsm_stall == 1'd0)) & (main_while_body_i_exitcond_reg == 1'd0))) */ begin
		main_while_body_i_indvar7 = main_while_body_i_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_1) & (fsm_stall == 1'd0))) begin
		main_while_body_i_indvar7_reg <= main_while_body_i_indvar7;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_body_i_4) & (fsm_stall == 1'd0)) & (main_while_body_i_exitcond_reg == 1'd0))) begin
		main_while_body_i_indvar7_reg <= main_while_body_i_indvar7;
	end
end
always @(*) begin
		main_while_body_i_dt_04_i = (1'd0 + (1 * {25'd0,main_while_body_i_indvar7_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_i_dt_04_i_reg <= main_while_body_i_dt_04_i;
	end
end
always @(*) begin
		main_while_body_i_st_05_i = (1'd0 + (1 * {25'd0,main_while_body_i_indvar7_reg}));
end
always @(*) begin
		main_while_body_i_0 = main_grid_out_a;
end
always @(*) begin
		main_while_body_i_1 = ({1'd0,main_while_body_i_indvar7_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_i_1_reg <= main_while_body_i_1;
	end
end
always @(*) begin
		main_while_body_i_exitcond = (main_while_body_i_1 == 32'd64);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_while_body_i_exitcond_reg <= main_while_body_i_exitcond;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i16_preheader_5) & (fsm_stall == 1'd0))) begin
		main_while_body_i16_indvar4 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_body_i16_8) & (fsm_stall == 1'd0)) & (main_while_body_i16_exitcond3_reg == 1'd0))) */ begin
		main_while_body_i16_indvar4 = main_while_body_i16_3_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i16_preheader_5) & (fsm_stall == 1'd0))) begin
		main_while_body_i16_indvar4_reg <= main_while_body_i16_indvar4;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_body_i16_8) & (fsm_stall == 1'd0)) & (main_while_body_i16_exitcond3_reg == 1'd0))) begin
		main_while_body_i16_indvar4_reg <= main_while_body_i16_indvar4;
	end
end
always @(*) begin
		main_while_body_i16_dt_05_i = (1'd0 + (4 * {27'd0,main_while_body_i16_indvar4_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_6)) begin
		main_while_body_i16_dt_05_i_reg <= main_while_body_i16_dt_05_i;
	end
end
always @(*) begin
		main_while_body_i16_st_06_i = (1'd0 + (4 * {27'd0,main_while_body_i16_indvar4_reg}));
end
always @(*) begin
		main_while_body_i16_2 = main_bypass_out_a;
end
always @(*) begin
		main_while_body_i16_3 = ({1'd0,main_while_body_i16_indvar4_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_6)) begin
		main_while_body_i16_3_reg <= main_while_body_i16_3;
	end
end
always @(*) begin
		main_while_body_i16_exitcond3 = (main_while_body_i16_3 == 32'd16);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_6)) begin
		main_while_body_i16_exitcond3_reg <= main_while_body_i16_exitcond3;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i10_preheader_9) & (fsm_stall == 1'd0))) begin
		main_while_body_i10_indvar1 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_body_i10_11) & (fsm_stall == 1'd0)) & (main_while_body_i10_exitcond2_reg == 1'd0))) */ begin
		main_while_body_i10_indvar1 = main_while_body_i10_4_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i10_preheader_9) & (fsm_stall == 1'd0))) begin
		main_while_body_i10_indvar1_reg <= main_while_body_i10_indvar1;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_body_i10_11) & (fsm_stall == 1'd0)) & (main_while_body_i10_exitcond2_reg == 1'd0))) begin
		main_while_body_i10_indvar1_reg <= main_while_body_i10_indvar1;
	end
end
always @(*) begin
		main_while_body_i10_s_010_i5 = (1'd0 + (4 * {29'd0,main_while_body_i10_indvar1_reg}));
end
always @(*) begin
		main_while_body_i10_4 = ({1'd0,main_while_body_i10_indvar1_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i10_10)) begin
		main_while_body_i10_4_reg <= main_while_body_i10_4;
	end
end
always @(*) begin
		main_while_body_i10_exitcond2 = (main_while_body_i10_4 == 32'd6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i10_10)) begin
		main_while_body_i10_exitcond2_reg <= main_while_body_i10_exitcond2;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i4_preheader_12) & (fsm_stall == 1'd0))) begin
		main_while_body_i4_indvar = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_while_body_i4_14) & (fsm_stall == 1'd0)) & (main_while_body_i4_exitcond1_reg == 1'd0))) */ begin
		main_while_body_i4_indvar = main_while_body_i4_5_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_while_body_i4_preheader_12) & (fsm_stall == 1'd0))) begin
		main_while_body_i4_indvar_reg <= main_while_body_i4_indvar;
	end
	if ((((cur_state == LEGUP_F_main_BB_while_body_i4_14) & (fsm_stall == 1'd0)) & (main_while_body_i4_exitcond1_reg == 1'd0))) begin
		main_while_body_i4_indvar_reg <= main_while_body_i4_indvar;
	end
end
always @(*) begin
		main_while_body_i4_s_010_i = (1'd0 + (4 * {29'd0,main_while_body_i4_indvar_reg}));
end
always @(*) begin
		main_while_body_i4_5 = ({1'd0,main_while_body_i4_indvar_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i4_13)) begin
		main_while_body_i4_5_reg <= main_while_body_i4_5;
	end
end
always @(*) begin
		main_while_body_i4_exitcond1 = (main_while_body_i4_5 == 32'd6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_while_body_i4_13)) begin
		main_while_body_i4_exitcond1_reg <= main_while_body_i4_exitcond1;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_state_0 = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_state_0 = main_sw_epilog_next_state_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_state_0_reg <= main_NodeBlock29_state_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_state_0_reg <= main_NodeBlock29_state_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_30_0 = 0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_current_sroa_30_0 = main_sw_epilog_next_current_sroa_6_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_30_0_reg <= main_NodeBlock29_current_sroa_30_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_30_0_reg <= main_NodeBlock29_current_sroa_30_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_0_0 = 0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_current_sroa_0_0 = main_sw_epilog_next_current_sroa_0_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_0_0_reg <= main_NodeBlock29_current_sroa_0_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_current_sroa_0_0_reg <= main_NodeBlock29_current_sroa_0_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_inputIndex_0 = 0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_inputIndex_0 = main_sw_epilog_next_inputIndex_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_inputIndex_0_reg <= main_NodeBlock29_inputIndex_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_inputIndex_0_reg <= main_NodeBlock29_inputIndex_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_stackIndex_0 = 0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_stackIndex_0 = main_sw_epilog_next_stackIndex_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_stackIndex_0_reg <= main_NodeBlock29_stackIndex_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_stackIndex_0_reg <= main_NodeBlock29_stackIndex_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_modified_0 = 1'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_modified_0 = main_sw_epilog_phitmp;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_modified_0_reg <= main_NodeBlock29_modified_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_modified_0_reg <= main_NodeBlock29_modified_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_firstEdge_0 = 1'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_firstEdge_0 = main_sw_epilog_phitmp279;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_firstEdge_0_reg <= main_NodeBlock29_firstEdge_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_firstEdge_0_reg <= main_NodeBlock29_firstEdge_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_state_0 = 0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_next_state_0 = main_sw_epilog_next_state_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_state_0_reg <= main_NodeBlock29_next_state_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_state_0_reg <= main_NodeBlock29_next_state_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_modified_0 = 8'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_next_modified_0 = main_sw_epilog_next_modified_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_modified_0_reg <= main_NodeBlock29_next_modified_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_modified_0_reg <= main_NodeBlock29_next_modified_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_firstEdge_0 = 8'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) */ begin
		main_NodeBlock29_next_firstEdge_0 = main_sw_epilog_next_firstEdge_1_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_NodeBlock29_preheader_15) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_firstEdge_0_reg <= main_NodeBlock29_next_firstEdge_0;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_epilog_98) & (fsm_stall == 1'd0))) begin
		main_NodeBlock29_next_firstEdge_0_reg <= main_NodeBlock29_next_firstEdge_0;
	end
end
always @(*) begin
		main_NodeBlock29_bit_select15 = main_NodeBlock29_current_sroa_30_0_reg[1:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock29_16)) begin
		main_NodeBlock29_bit_select15_reg <= main_NodeBlock29_bit_select15;
	end
end
always @(*) begin
		main_NodeBlock29_bit_select13 = main_NodeBlock29_current_sroa_0_0_reg[1:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock29_16)) begin
		main_NodeBlock29_bit_select13_reg <= main_NodeBlock29_bit_select13;
	end
end
always @(*) begin
		main_NodeBlock29_bit_select11 = main_NodeBlock29_current_sroa_30_0_reg[31:2];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock29_16)) begin
		main_NodeBlock29_bit_select11_reg <= main_NodeBlock29_bit_select11;
	end
end
always @(*) begin
		main_NodeBlock29_bit_select9 = main_NodeBlock29_current_sroa_0_0_reg[31:2];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock29_16)) begin
		main_NodeBlock29_bit_select9_reg <= main_NodeBlock29_bit_select9;
	end
end
always @(*) begin
		main_NodeBlock29_bit_select5 = main_NodeBlock29_current_sroa_0_0_reg[29:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock29_16)) begin
		main_NodeBlock29_bit_select5_reg <= main_NodeBlock29_bit_select5;
	end
end
always @(*) begin
		main_NodeBlock29_Pivot30 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock29_Pivot30_op1_temp}));
end
always @(*) begin
		main_NodeBlock27_Pivot28 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock27_Pivot28_op1_temp}));
end
always @(*) begin
		main_NodeBlock25_Pivot26 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock25_Pivot26_op1_temp}));
end
always @(*) begin
		main_NodeBlock23_Pivot24 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock23_Pivot24_op1_temp}));
end
always @(*) begin
		main_LeafBlock21_SwitchLeaf22 = (main_NodeBlock29_state_0_reg == 32'd15);
end
always @(*) begin
		main_NodeBlock19_Pivot20 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock19_Pivot20_op1_temp}));
end
always @(*) begin
		main_NodeBlock17_Pivot18 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock17_Pivot18_op1_temp}));
end
always @(*) begin
		main_NodeBlock15_Pivot16 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock15_Pivot16_op1_temp}));
end
always @(*) begin
		main_NodeBlock15_bit_concat23 = {main_NodeBlock29_bit_select5_reg[29:0], main_NodeBlock15_bit_concat23_bit_select_operand_2[1:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock15_23)) begin
		main_NodeBlock15_bit_concat23_reg <= main_NodeBlock15_bit_concat23;
	end
end
always @(*) begin
		main_NodeBlock13_Pivot14 = ($signed(main_NodeBlock29_state_0_reg) < $signed({26'd0,main_NodeBlock13_Pivot14_op1_temp}));
end
always @(*) begin
		main_NodeBlock11_Pivot12 = ($signed(main_NodeBlock29_state_0_reg) < $signed({27'd0,main_NodeBlock11_Pivot12_op1_temp}));
end
always @(*) begin
		main_NodeBlock9_Pivot10 = ($signed(main_NodeBlock29_state_0_reg) < $signed({27'd0,main_NodeBlock9_Pivot10_op1_temp}));
end
always @(*) begin
		main_NodeBlock7_Pivot8 = ($signed(main_NodeBlock29_state_0_reg) < $signed({27'd0,main_NodeBlock7_Pivot8_op1_temp}));
end
always @(*) begin
		main_NodeBlock7_bit_concat22 = {main_NodeBlock29_bit_select5_reg[29:0], main_NodeBlock7_bit_concat22_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_NodeBlock7_arrayidx32 = (1'd0 + (1 * main_NodeBlock7_bit_concat22));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock7_27)) begin
		main_NodeBlock7_arrayidx32_reg <= main_NodeBlock7_arrayidx32;
	end
end
always @(*) begin
		main_NodeBlock5_Pivot6 = ($signed(main_NodeBlock29_state_0_reg) < $signed({27'd0,main_NodeBlock5_Pivot6_op1_temp}));
end
always @(*) begin
		main_NodeBlock5_bit_concat21 = {main_NodeBlock29_bit_select5_reg[29:0], main_NodeBlock5_bit_concat21_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_NodeBlock5_arrayidx62 = (1'd0 + (1 * main_NodeBlock5_bit_concat21));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_NodeBlock5_28)) begin
		main_NodeBlock5_arrayidx62_reg <= main_NodeBlock5_arrayidx62;
	end
end
always @(*) begin
		main_NodeBlock3_Pivot4 = ($signed(main_NodeBlock29_state_0_reg) < $signed({28'd0,main_NodeBlock3_Pivot4_op1_temp}));
end
always @(*) begin
		main_NodeBlock1_Pivot2 = ($signed(main_NodeBlock29_state_0_reg) < $signed({28'd0,main_NodeBlock1_Pivot2_op1_temp}));
end
always @(*) begin
		main_NodeBlock_Pivot = ($signed(main_NodeBlock29_state_0_reg) < $signed({29'd0,main_NodeBlock_Pivot_op1_temp}));
end
always @(*) begin
		main_LeafBlock_SwitchLeaf = (main_NodeBlock29_state_0_reg == 32'd0);
end
always @(*) begin
		main_sw_bb1_arrayidx = (1'd0 + (4 * main_NodeBlock29_inputIndex_0_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb1_33)) begin
		main_sw_bb1_arrayidx_reg <= main_sw_bb1_arrayidx;
	end
end
always @(*) begin
		main_sw_bb1_6 = (32'd49157 >>> (main_NodeBlock29_inputIndex_0_reg % 32));
end
always @(*) begin
		main_sw_bb1_bit_select19 = main_sw_bb1_6[0];
end
always @(*) begin
		main_sw_bb1_bit_concat20 = {main_sw_bb1_bit_concat20_bit_select_operand_0[30:0], main_sw_bb1_bit_select19};
end
always @(*) begin
		main_sw_bb1_cmp = (main_sw_bb1_bit_concat20 == 32'd0);
end
always @(*) begin
		main_sw_bb1_add8_pre = (main_NodeBlock29_inputIndex_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb1_33)) begin
		main_sw_bb1_add8_pre_reg <= main_sw_bb1_add8_pre;
	end
end
always @(*) begin
		main_land_lhs_true_7 = (32'd49157 >>> (main_sw_bb1_add8_pre_reg % 32));
end
always @(*) begin
		main_land_lhs_true_bit_select17 = main_land_lhs_true_7[0];
end
always @(*) begin
		main_land_lhs_true_bit_concat18 = {main_land_lhs_true_bit_concat18_bit_select_operand_0[30:0], main_land_lhs_true_bit_select17};
end
always @(*) begin
		main_land_lhs_true_cmp4 = (main_land_lhs_true_bit_concat18 == 32'd0);
end
always @(*) begin
		main_if_else_8 = main_input_out_a;
end
always @(*) begin
		main_if_else_arrayidx9 = (1'd0 + (4 * main_sw_bb1_add8_pre_reg));
end
always @(*) begin
		main_if_else_9 = main_input_out_b;
end
always @(*) begin
		main_if_else_add11 = (main_NodeBlock29_inputIndex_0_reg + 32'd2);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_else_35)) begin
		main_if_else_add11_reg <= main_if_else_add11;
	end
end
always @(*) begin
		main_sw_bb12_bit_concat16 = {main_sw_bb12_bit_concat16_bit_select_operand_0[29:0], main_NodeBlock29_bit_select15_reg[1:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb12_37)) begin
		main_sw_bb12_bit_concat16_reg <= main_sw_bb12_bit_concat16;
	end
end
always @(*) begin
		main_sw_bb12_bit_concat14 = {main_sw_bb12_bit_concat14_bit_select_operand_0[29:0], main_NodeBlock29_bit_select13_reg[1:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb12_37)) begin
		main_sw_bb12_bit_concat14_reg <= main_sw_bb12_bit_concat14;
	end
end
always @(*) begin
		main_sw_bb12_cmp16 = (main_sw_bb12_bit_concat16 == main_sw_bb12_bit_concat14);
end
always @(*) begin
		main_if_else18_sub = (main_sw_bb12_bit_concat16_reg - main_sw_bb12_bit_concat14_reg);
end
always @(*) begin
		main_if_else18_cmp24 = ($signed(main_if_else18_sub) > $signed({30'd0,main_if_else18_cmp24_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_else18_38)) begin
		main_if_else18_cmp24_reg <= main_if_else18_cmp24;
	end
end
always @(*) begin
		main_if_else18_1 = (main_if_else18_cmp24_reg ? 32'd6 : 32'd4);
end
always @(*) begin
		main_sw_bb29_10 = main_entry_grid_out_a;
end
always @(*) begin
		main_sw_bb29_tobool = (main_sw_bb29_10 == 8'd0);
end
always @(*) begin
		main_lor_lhs_false_arrayidx34 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(*) begin
		main_lor_lhs_false_11 = main_entry_bypass_out_a;
end
always @(*) begin
		main_lor_lhs_false_cmp35_not = (main_lor_lhs_false_11 < 32'd2);
end
always @(*) begin
		main_lor_lhs_false_brmerge = (main_lor_lhs_false_cmp35_not | main_NodeBlock29_firstEdge_0_reg);
end
always @(*) begin
		main_lor_lhs_false_292 = (main_lor_lhs_false_brmerge ? 32'd7 : 32'd8);
end
always @(*) begin
		main_if_then47_arrayidx49 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then47_46)) begin
		main_if_then47_arrayidx49_reg <= main_if_then47_arrayidx49;
	end
end
always @(*) begin
		main_if_then47_12 = main_entry_bypass_out_a;
end
always @(*) begin
		main_if_then47_inc = (main_if_then47_12 + 32'd1);
end
always @(*) begin
		main_if_end50_add52 = (main_NodeBlock29_current_sroa_0_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_if_end50_add52_reg <= main_if_end50_add52;
	end
end
always @(*) begin
		main_if_end50_arrayidx55 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end50_arrayidx56 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end50_add57 = (main_NodeBlock29_stackIndex_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_if_end50_add57_reg <= main_if_end50_add57;
	end
end
always @(*) begin
		main_sw_bb58_13 = main_entry_grid_out_a;
end
always @(*) begin
		main_sw_bb58_tobool63 = (main_sw_bb58_13 == 8'd0);
end
always @(*) begin
		main_lor_lhs_false64_arrayidx66 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(*) begin
		main_lor_lhs_false64_14 = main_entry_bypass_out_a;
end
always @(*) begin
		main_lor_lhs_false64_cmp67_not = (main_lor_lhs_false64_14 < 32'd3);
end
always @(*) begin
		main_lor_lhs_false64_brmerge286 = (main_lor_lhs_false64_cmp67_not | main_NodeBlock29_firstEdge_0_reg);
end
always @(*) begin
		main_lor_lhs_false64_293 = (main_lor_lhs_false64_brmerge286 ? 32'd5 : 32'd8);
end
always @(*) begin
		main_if_then79_arrayidx81 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then79_57)) begin
		main_if_then79_arrayidx81_reg <= main_if_then79_arrayidx81;
	end
end
always @(*) begin
		main_if_then79_15 = main_entry_bypass_out_a;
end
always @(*) begin
		main_if_then79_inc82 = (main_if_then79_15 + 32'd1);
end
always @(*) begin
		main_if_end83_sub85 = (main_NodeBlock29_current_sroa_0_0_reg + $signed(-32'd1));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_if_end83_sub85_reg <= main_if_end83_sub85;
	end
end
always @(*) begin
		main_if_end83_arrayidx88 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end83_arrayidx89 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end83_add90 = (main_NodeBlock29_stackIndex_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_if_end83_add90_reg <= main_if_end83_add90;
	end
end
always @(*) begin
		main_sw_bb91_bit_concat12 = {main_sw_bb91_bit_concat12_bit_select_operand_0[1:0], main_NodeBlock29_bit_select11_reg[29:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb91_62)) begin
		main_sw_bb91_bit_concat12_reg <= main_sw_bb91_bit_concat12;
	end
end
always @(*) begin
		main_sw_bb91_bit_concat10 = {main_sw_bb91_bit_concat10_bit_select_operand_0[1:0], main_NodeBlock29_bit_select9_reg[29:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb91_62)) begin
		main_sw_bb91_bit_concat10_reg <= main_sw_bb91_bit_concat10;
	end
end
always @(*) begin
		main_sw_bb91_cmp96 = (main_sw_bb91_bit_concat12 == main_sw_bb91_bit_concat10);
end
always @(*) begin
		main_if_else98_sub95 = (main_sw_bb91_bit_concat12_reg - main_sw_bb91_bit_concat10_reg);
end
always @(*) begin
		main_if_else98_cmp104 = ($signed(main_if_else98_sub95) > $signed({30'd0,main_if_else98_cmp104_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_else98_63)) begin
		main_if_else98_cmp104_reg <= main_if_else98_cmp104;
	end
end
always @(*) begin
		main_if_else98_287 = (main_if_else98_cmp104_reg ? 32'd11 : 32'd9);
end
always @(*) begin
		main_sw_bb109_bit_concat8 = {main_NodeBlock29_bit_select5_reg[29:0], main_sw_bb109_bit_concat8_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_sw_bb109_arrayidx113 = (1'd0 + (1 * main_sw_bb109_bit_concat8));
end
always @(*) begin
		main_sw_bb109_16 = main_entry_grid_out_a;
end
always @(*) begin
		main_sw_bb109_tobool114 = (main_sw_bb109_16 == 8'd0);
end
always @(*) begin
		main_lor_lhs_false115_arrayidx117 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(*) begin
		main_lor_lhs_false115_17 = main_entry_bypass_out_a;
end
always @(*) begin
		main_lor_lhs_false115_cmp118_not = (main_lor_lhs_false115_17 < 32'd2);
end
always @(*) begin
		main_lor_lhs_false115_brmerge288 = (main_lor_lhs_false115_cmp118_not | main_NodeBlock29_firstEdge_0_reg);
end
always @(*) begin
		main_lor_lhs_false115_294 = (main_lor_lhs_false115_brmerge288 ? 32'd12 : 32'd13);
end
always @(*) begin
		main_sw_bb124_bit_concat7 = {main_NodeBlock29_bit_select5_reg[29:0], main_sw_bb124_bit_concat7_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_sw_bb124_arrayidx128 = (1'd0 + (1 * main_sw_bb124_bit_concat7));
end
always @(*) begin
		main_if_then130_arrayidx132 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then130_71)) begin
		main_if_then130_arrayidx132_reg <= main_if_then130_arrayidx132;
	end
end
always @(*) begin
		main_if_then130_18 = main_entry_bypass_out_a;
end
always @(*) begin
		main_if_then130_inc133 = (main_if_then130_18 + 32'd1);
end
always @(*) begin
		main_if_end134_add136 = (main_NodeBlock29_current_sroa_0_0_reg + 32'd4);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_if_end134_add136_reg <= main_if_end134_add136;
	end
end
always @(*) begin
		main_if_end134_arrayidx139 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end134_arrayidx140 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end134_add141 = (main_NodeBlock29_stackIndex_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_if_end134_add141_reg <= main_if_end134_add141;
	end
end
always @(*) begin
		main_sw_bb142_bit_concat6 = {main_NodeBlock29_bit_select5_reg[29:0], main_sw_bb142_bit_concat6_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_sw_bb142_arrayidx146 = (1'd0 + (1 * main_sw_bb142_bit_concat6));
end
always @(*) begin
		main_sw_bb142_19 = main_entry_grid_out_a;
end
always @(*) begin
		main_sw_bb142_tobool147 = (main_sw_bb142_19 == 8'd0);
end
always @(*) begin
		main_lor_lhs_false148_arrayidx150 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(*) begin
		main_lor_lhs_false148_20 = main_entry_bypass_out_a;
end
always @(*) begin
		main_lor_lhs_false148_cmp151_not = (main_lor_lhs_false148_20 < 32'd3);
end
always @(*) begin
		main_lor_lhs_false148_brmerge289 = (main_lor_lhs_false148_cmp151_not | main_NodeBlock29_firstEdge_0_reg);
end
always @(*) begin
		main_lor_lhs_false148_295 = (main_lor_lhs_false148_brmerge289 ? 32'd10 : 32'd13);
end
always @(*) begin
		main_sw_bb157_arrayidx161 = (1'd0 + (1 * main_NodeBlock15_bit_concat23_reg));
end
always @(*) begin
		main_if_then163_arrayidx165 = (1'd0 + (4 * main_NodeBlock29_current_sroa_0_0_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then163_82)) begin
		main_if_then163_arrayidx165_reg <= main_if_then163_arrayidx165;
	end
end
always @(*) begin
		main_if_then163_21 = main_entry_bypass_out_a;
end
always @(*) begin
		main_if_then163_inc166 = (main_if_then163_21 + 32'd1);
end
always @(*) begin
		main_if_end167_sub169 = (main_NodeBlock29_current_sroa_0_0_reg + $signed(-32'd4));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_if_end167_sub169_reg <= main_if_end167_sub169;
	end
end
always @(*) begin
		main_if_end167_arrayidx172 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end167_arrayidx173 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_if_end167_add174 = (main_NodeBlock29_stackIndex_0_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_if_end167_add174_reg <= main_if_end167_add174;
	end
end
always @(*) begin
		main_sw_bb175_cmp178 = (main_NodeBlock29_current_sroa_0_0_reg == main_NodeBlock29_current_sroa_30_0_reg);
end
always @(*) begin
		main_sw_bb175_290 = (main_sw_bb175_cmp178 ? 32'd1 : 32'd14);
end
always @(*) begin
		main_sw_bb182_291 = (main_NodeBlock29_modified_0_reg ? 32'd3 : 32'd15);
end
always @(*) begin
		main_sw_bb182_next_modified_0 = (main_NodeBlock29_modified_0_reg ? 8'd0 : main_NodeBlock29_next_modified_0_reg);
end
always @(*) begin
		main_sw_bb187_arrayidx188 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_sw_bb187_22 = main_entry_stackNode_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_90)) begin
		main_sw_bb187_22_reg <= main_sw_bb187_22;
	end
end
always @(*) begin
		main_sw_bb187_bit_select3 = main_sw_bb187_22[29:0];
end
always @(*) begin
		main_sw_bb187_bit_concat4 = {main_sw_bb187_bit_select3[29:0], main_sw_bb187_bit_concat4_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_sw_bb187_arrayidx190 = (1'd0 + (4 * main_NodeBlock29_stackIndex_0_reg));
end
always @(*) begin
		main_sw_bb187_23 = main_entry_stackOutput_out_a;
end
always @(*) begin
		main_sw_bb187_add191 = (main_sw_bb187_bit_concat4 + main_sw_bb187_23);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_90)) begin
		main_sw_bb187_add191_reg <= main_sw_bb187_add191;
	end
end
always @(*) begin
		main_sw_bb187_arrayidx192 = (1'd0 + (1 * main_sw_bb187_add191_reg));
end
always @(*) begin
		main_sw_bb187_cmp193 = (main_NodeBlock29_stackIndex_0_reg == 32'd0);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_89)) begin
		main_sw_bb187_cmp193_reg <= main_sw_bb187_cmp193;
	end
end
always @(*) begin
		main_if_else195_sub196 = (main_NodeBlock29_stackIndex_0_reg + $signed(-32'd1));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_else195_93)) begin
		main_if_else195_sub196_reg <= main_if_else195_sub196;
	end
end
always @(*) begin
		main_if_else195_arrayidx198 = (1'd0 + (4 * main_sw_bb187_22_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_else195_93)) begin
		main_if_else195_arrayidx198_reg <= main_if_else195_arrayidx198;
	end
end
always @(*) begin
		main_if_else195_24 = main_entry_bypass_out_a;
end
always @(*) begin
		main_if_else195_dec = (main_if_else195_24 + $signed(-32'd1));
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_state_1 = 32'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd2;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd3;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_state_1 = 32'd8;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {29'd0,main_if_else18_1};
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd8;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_lor_lhs_false_292};
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd3;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd8;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_lor_lhs_false64_293};
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd3;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_state_1 = 32'd13;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_if_else98_287};
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd13;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_lor_lhs_false115_294};
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd8;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd13;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_lor_lhs_false148_295};
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd8;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_sw_bb175_290};
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = {28'd0,main_sw_bb182_291};
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_state_1 = 32'd1;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1 = 32'd15;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_state_1 = main_NodeBlock29_next_state_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_state_1_reg <= main_sw_epilog_next_state_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_if_else_9;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_current_sroa_6_1 = main_NodeBlock29_current_sroa_30_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_6_1_reg <= main_sw_epilog_next_current_sroa_6_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_if_else_8;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_if_end50_add52_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_if_end83_sub85_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_if_end134_add136_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_if_end167_sub169_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_current_sroa_0_1 = main_NodeBlock29_current_sroa_0_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_current_sroa_0_1_reg <= main_sw_epilog_next_current_sroa_0_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_if_else_add11_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_inputIndex_1 = main_NodeBlock29_inputIndex_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_inputIndex_1_reg <= main_sw_epilog_next_inputIndex_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = 32'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_if_end50_add57_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_if_end83_add90_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_if_end134_add141_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_if_end167_add174_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1 = 32'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1 = main_if_else195_sub196_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_stackIndex_1 = main_NodeBlock29_stackIndex_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_stackIndex_1_reg <= main_sw_epilog_next_stackIndex_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = 8'd1;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_sw_bb182_next_modified_0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_modified_1 = main_NodeBlock29_next_modified_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_modified_1_reg <= main_sw_epilog_next_modified_1;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = 8'd1;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = 8'd0;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = 8'd0;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) */ begin
		main_sw_epilog_next_firstEdge_1 = main_NodeBlock29_next_firstEdge_0_reg;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_32) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_land_lhs_true_34) & (fsm_stall == 1'd0)) & (main_land_lhs_true_cmp4 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else_36) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb12_37) & (fsm_stall == 1'd0)) & (main_sw_bb12_cmp16 == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else18_39) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb29_41) & (fsm_stall == 1'd0)) & (main_sw_bb29_tobool == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false_43) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end50_50) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb58_52) & (fsm_stall == 1'd0)) & (main_sw_bb58_tobool63 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false64_54) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end83_61) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb91_62) & (fsm_stall == 1'd0)) & (main_sw_bb91_cmp96 == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else98_64) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb109_66) & (fsm_stall == 1'd0)) & (main_sw_bb109_tobool114 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false115_68) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end134_75) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb142_77) & (fsm_stall == 1'd0)) & (main_sw_bb142_tobool147 == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_lor_lhs_false148_79) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_end167_86) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb175_87) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_sw_bb182_88) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_sw_bb187_92) & (fsm_stall == 1'd0)) & (main_sw_bb187_cmp193_reg == 1'd1))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_if_else195_95) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
	if (((cur_state == LEGUP_F_main_BB_NewDefault_97) & (fsm_stall == 1'd0))) begin
		main_sw_epilog_next_firstEdge_1_reg <= main_sw_epilog_next_firstEdge_1;
	end
end
always @(*) begin
		main_sw_epilog_bit_select1 = main_sw_epilog_next_modified_1_reg[0];
end
always @(*) begin
		main_sw_epilog_bit_select = main_sw_epilog_next_firstEdge_1_reg[0];
end
always @(*) begin
		main_sw_epilog_bit_concat2 = {main_sw_epilog_bit_concat2_bit_select_operand_0[6:0], main_sw_epilog_bit_select1};
end
always @(*) begin
		main_sw_epilog_phitmp = (main_sw_epilog_bit_concat2 != 8'd0);
end
always @(*) begin
		main_sw_epilog_bit_concat = {main_sw_epilog_bit_concat_bit_select_operand_0[6:0], main_sw_epilog_bit_select};
end
always @(*) begin
		main_sw_epilog_phitmp279 = (main_sw_epilog_bit_concat != 8'd0);
end
always @(*) begin
	main_input_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_else_35)) begin
		main_input_address_a = (main_sw_bb1_arrayidx_reg >>> 3'd2);
	end
end
always @(*) begin
	main_input_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_else_35)) begin
		main_input_address_b = (main_if_else_arrayidx9 >>> 3'd2);
	end
end
always @(*) begin
	main_grid_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_2)) begin
		main_grid_address_a = (main_while_body_i_st_05_i >>> 3'd0);
	end
end
assign main_grid_address_b = 'dx;
always @(*) begin
	main_bypass_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_6)) begin
		main_bypass_address_a = (main_while_body_i16_st_06_i >>> 3'd2);
	end
end
assign main_bypass_address_b = 'dx;
always @(*) begin
	main_entry_grid_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_3)) begin
		main_entry_grid_address_a = (main_while_body_i_dt_04_i_reg >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb29_40)) begin
		main_entry_grid_address_a = (main_NodeBlock7_arrayidx32_reg >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb41_44)) begin
		main_entry_grid_address_a = (main_NodeBlock7_arrayidx32_reg >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb58_51)) begin
		main_entry_grid_address_a = (main_NodeBlock5_arrayidx62_reg >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb73_55)) begin
		main_entry_grid_address_a = (main_NodeBlock5_arrayidx62_reg >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb109_65)) begin
		main_entry_grid_address_a = (main_sw_bb109_arrayidx113 >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb124_69)) begin
		main_entry_grid_address_a = (main_sw_bb124_arrayidx128 >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb142_76)) begin
		main_entry_grid_address_a = (main_sw_bb142_arrayidx146 >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb157_80)) begin
		main_entry_grid_address_a = (main_sw_bb157_arrayidx161 >>> 3'd0);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_91)) begin
		main_entry_grid_address_a = (main_sw_bb187_arrayidx192 >>> 3'd0);
	end
end
always @(*) begin
	main_entry_grid_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_3)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb41_44)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb73_55)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb124_69)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb157_80)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_91)) begin
		main_entry_grid_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_grid_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i_3)) begin
		main_entry_grid_in_a = main_while_body_i_0;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb41_44)) begin
		main_entry_grid_in_a = 8'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb73_55)) begin
		main_entry_grid_in_a = 8'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb124_69)) begin
		main_entry_grid_in_a = 8'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb157_80)) begin
		main_entry_grid_in_a = 8'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_91)) begin
		main_entry_grid_in_a = 8'd0;
	end
end
always @(*) begin
	main_entry_bypass_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_7)) begin
		main_entry_bypass_address_a = (main_while_body_i16_dt_05_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_lor_lhs_false_42)) begin
		main_entry_bypass_address_a = (main_lor_lhs_false_arrayidx34 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_46)) begin
		main_entry_bypass_address_a = (main_if_then47_arrayidx49 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_47)) begin
		main_entry_bypass_address_a = (main_if_then47_arrayidx49_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_lor_lhs_false64_53)) begin
		main_entry_bypass_address_a = (main_lor_lhs_false64_arrayidx66 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then79_57)) begin
		main_entry_bypass_address_a = (main_if_then79_arrayidx81 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then79_58)) begin
		main_entry_bypass_address_a = (main_if_then79_arrayidx81_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_lor_lhs_false115_67)) begin
		main_entry_bypass_address_a = (main_lor_lhs_false115_arrayidx117 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then130_71)) begin
		main_entry_bypass_address_a = (main_if_then130_arrayidx132 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then130_72)) begin
		main_entry_bypass_address_a = (main_if_then130_arrayidx132_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_lor_lhs_false148_78)) begin
		main_entry_bypass_address_a = (main_lor_lhs_false148_arrayidx150 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then163_82)) begin
		main_entry_bypass_address_a = (main_if_then163_arrayidx165 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then163_83)) begin
		main_entry_bypass_address_a = (main_if_then163_arrayidx165_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_else195_93)) begin
		main_entry_bypass_address_a = (main_if_else195_arrayidx198 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_else195_94)) begin
		main_entry_bypass_address_a = (main_if_else195_arrayidx198_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_bypass_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_7)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_47)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then79_58)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then130_72)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then163_83)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_else195_94)) begin
		main_entry_bypass_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_bypass_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i16_7)) begin
		main_entry_bypass_in_a = main_while_body_i16_2;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then47_47)) begin
		main_entry_bypass_in_a = main_if_then47_inc;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then79_58)) begin
		main_entry_bypass_in_a = main_if_then79_inc82;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then130_72)) begin
		main_entry_bypass_in_a = main_if_then130_inc133;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then163_83)) begin
		main_entry_bypass_in_a = main_if_then163_inc166;
	end
	if ((cur_state == LEGUP_F_main_BB_if_else195_94)) begin
		main_entry_bypass_in_a = main_if_else195_dec;
	end
end
always @(*) begin
	main_entry_stackNode_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i10_10)) begin
		main_entry_stackNode_address_a = (main_while_body_i10_s_010_i5 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackNode_address_a = (main_if_end50_arrayidx55 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackNode_address_a = (main_if_end83_arrayidx88 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackNode_address_a = (main_if_end134_arrayidx139 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackNode_address_a = (main_if_end167_arrayidx172 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_89)) begin
		main_entry_stackNode_address_a = (main_sw_bb187_arrayidx188 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_stackNode_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_while_body_i10_10)) begin
		main_entry_stackNode_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackNode_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackNode_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackNode_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackNode_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_stackNode_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i10_10)) begin
		main_entry_stackNode_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackNode_in_a = main_NodeBlock29_current_sroa_0_0_reg;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackNode_in_a = main_NodeBlock29_current_sroa_0_0_reg;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackNode_in_a = main_NodeBlock29_current_sroa_0_0_reg;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackNode_in_a = main_NodeBlock29_current_sroa_0_0_reg;
	end
end
always @(*) begin
	main_entry_stackOutput_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i4_13)) begin
		main_entry_stackOutput_address_a = (main_while_body_i4_s_010_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackOutput_address_a = (main_if_end50_arrayidx56 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackOutput_address_a = (main_if_end83_arrayidx89 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackOutput_address_a = (main_if_end134_arrayidx140 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackOutput_address_a = (main_if_end167_arrayidx173 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb187_89)) begin
		main_entry_stackOutput_address_a = (main_sw_bb187_arrayidx190 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_stackOutput_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_while_body_i4_13)) begin
		main_entry_stackOutput_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackOutput_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackOutput_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackOutput_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackOutput_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_stackOutput_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_while_body_i4_13)) begin
		main_entry_stackOutput_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end50_49)) begin
		main_entry_stackOutput_in_a = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end83_60)) begin
		main_entry_stackOutput_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end134_74)) begin
		main_entry_stackOutput_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_end167_85)) begin
		main_entry_stackOutput_in_a = 32'd0;
	end
end
assign main_NodeBlock29_Pivot30_op1_temp = 32'd8;
assign main_NodeBlock27_Pivot28_op1_temp = 32'd12;
assign main_NodeBlock25_Pivot26_op1_temp = 32'd14;
assign main_NodeBlock23_Pivot24_op1_temp = 32'd15;
assign main_NodeBlock19_Pivot20_op1_temp = 32'd13;
assign main_NodeBlock17_Pivot18_op1_temp = 32'd10;
assign main_NodeBlock15_Pivot16_op1_temp = 32'd11;
assign main_NodeBlock15_bit_concat23_bit_select_operand_2 = 2'd0;
assign main_NodeBlock13_Pivot14_op1_temp = 32'd9;
assign main_NodeBlock11_Pivot12_op1_temp = 32'd4;
assign main_NodeBlock9_Pivot10_op1_temp = 32'd6;
assign main_NodeBlock7_Pivot8_op1_temp = 32'd7;
assign main_NodeBlock7_bit_concat22_bit_select_operand_2 = -2'd1;
assign main_NodeBlock5_Pivot6_op1_temp = 32'd5;
assign main_NodeBlock5_bit_concat21_bit_select_operand_2 = -2'd2;
assign main_NodeBlock3_Pivot4_op1_temp = 32'd2;
assign main_NodeBlock1_Pivot2_op1_temp = 32'd3;
assign main_NodeBlock_Pivot_op1_temp = 32'd1;
assign main_sw_bb1_bit_concat20_bit_select_operand_0 = 31'd0;
assign main_land_lhs_true_bit_concat18_bit_select_operand_0 = 31'd0;
assign main_sw_bb12_bit_concat16_bit_select_operand_0 = 30'd0;
assign main_sw_bb12_bit_concat14_bit_select_operand_0 = 30'd0;
assign main_if_else18_cmp24_op1_temp = 32'd0;
assign main_sw_bb91_bit_concat12_bit_select_operand_0 = 2'd0;
assign main_sw_bb91_bit_concat10_bit_select_operand_0 = 2'd0;
assign main_if_else98_cmp104_op1_temp = 32'd0;
assign main_sw_bb109_bit_concat8_bit_select_operand_2 = 2'd1;
assign main_sw_bb124_bit_concat7_bit_select_operand_2 = 2'd1;
assign main_sw_bb142_bit_concat6_bit_select_operand_2 = 2'd0;
assign main_sw_bb187_bit_concat4_bit_select_operand_2 = 2'd0;
assign main_sw_epilog_bit_concat2_bit_select_operand_0 = 7'd0;
assign main_sw_epilog_bit_concat_bit_select_operand_0 = 7'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb200_96)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_sw_bb200_96)) begin
		return_val <= 32'd1;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module rom_dual_port
(
	clk,
	clken,
	address_a,
	q_a,
	address_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  init_file = {`MEM_INIT_DIR, "UNUSED.mif"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;

(* ram_init_file = init_file *) reg [width_a-1:0] ram [numwords_a-1:0];

integer i;
/* synthesis translate_off */
ALTERA_MF_MEMORY_INITIALIZATION mem ();
reg [8*256:1] ram_ver_file;
initial begin
	if (init_file == {`MEM_INIT_DIR, "UNUSED.mif"})
    begin
		for (i = 0; i < numwords_a; i = i + 1)
			ram[i] = 0;
    end
	else
    begin
        // modelsim can't read .mif files directly. So use Altera function to
        // convert them to .ver files
        mem.convert_to_ver_file(init_file, width_a, ram_ver_file);
        $readmemh(ram_ver_file, ram);
    end
end
/* synthesis translate_on */

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  address_b_reg[0] = address_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
   end
end

always @ (posedge clk)
if (clken)
begin
    q_a_wire <= ram[address_a_reg[input_latency]];
end

always @ (posedge clk)
if (clken)
begin
    q_b_wire <= ram[address_b_reg[input_latency]];
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
